`include "CPU.vh"

// Asynchronous ROM (Program Memory)

module AsyncROM(
	// You fill this in...
);


endmodule

